`timescale 1ns/1ps
// Name: mux32_8x1_tb.v
// Module: MUX32_8x1_TB
// Input: 
// Output: 
//
// Notes: Common definitions
// 
//
// Revision History:
//
// Version	Date		Who		email			note
//------------------------------------------------------------------------------------------
//  1.0     Apr 18, 2020	Ryan Tran	tranryanp@gmail.com	Initial creation
//------------------------------------------------------------------------------------------

module MUX32_8x1_TB;
reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7;
reg [2:0] S;
wire [31:0] Y;

MUX32_8x1 mux32_8x1_inst1(.Y(Y), .I0(I0), .I1(I1), .I2(I2), .I3(I3),
			  .I4(I4), .I5(I5), .I6(I6), .I7(I7), .S(S));

initial
begin
I0 = 0; I1 = 0; I2 = 0; I3 = 0; I4 = 0; I5 = 0; I6 = 0; I7 = 0; S = 0;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, S:%d Y:%d\n",
I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703;
I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; S = 0;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, S:%d Y:%d\n",
I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703;
I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; S = 1;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, S:%d Y:%d\n",
I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703;
I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; S = 2;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, S:%d Y:%d\n",
I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703;
I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; S = 3;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, S:%d Y:%d\n",
I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703;
I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; S = 4;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, S:%d Y:%d\n",
I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703;
I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; S = 5;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, S:%d Y:%d\n",
I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703;
I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; S = 6;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, S:%d Y:%d\n",
I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703;
I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; S = 7;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, S:%d Y:%d\n",
I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
end

endmodule
