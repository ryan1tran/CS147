`timescale 1ns/1ps

module MUX32_8x1_TB;
wire [31:0] Y;
reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7;
reg [2:0] S;

MUX32_8x1 mux32_8x1_inst(.Y(Y), .I0(I0), .I1(I1), .I2(I2), .I3(I3),
                         .I4(I4), .I5(I5), .I6(I6), .I7(I7), .S(S));

initial
begin
I0 = 0; I1 = 0; I2 = 0; I3 = 0; I4 = 0; I5 = 0; I6 = 0; I7 = 0; S = 0;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
#5 I0 = 4294967288; I1 = 4294967289; I2 = 4294967290; I3 = 4294967291; I4 = 4294967292; I5 = 4294967293; I6 = 4294967294; I7 = 4294967295; S = 0;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
#5 I0 = 4294967288; I1 = 4294967289; I2 = 4294967290; I3 = 4294967291; I4 = 4294967292; I5 = 4294967293; I6 = 4294967294; I7 = 4294967295; S = 1;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
#5 I0 = 4294967288; I1 = 4294967289; I2 = 4294967290; I3 = 4294967291; I4 = 4294967292; I5 = 4294967293; I6 = 4294967294; I7 = 4294967295; S = 2;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
#5 I0 = 4294967288; I1 = 4294967289; I2 = 4294967290; I3 = 4294967291; I4 = 4294967292; I5 = 4294967293; I6 = 4294967294; I7 = 4294967295; S = 3;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
#5 I0 = 4294967288; I1 = 4294967289; I2 = 4294967290; I3 = 4294967291; I4 = 4294967292; I5 = 4294967293; I6 = 4294967294; I7 = 4294967295; S = 4;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
#5 I0 = 4294967288; I1 = 4294967289; I2 = 4294967290; I3 = 4294967291; I4 = 4294967292; I5 = 4294967293; I6 = 4294967294; I7 = 4294967295; S = 5;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
#5 I0 = 4294967288; I1 = 4294967289; I2 = 4294967290; I3 = 4294967291; I4 = 4294967292; I5 = 4294967293; I6 = 4294967294; I7 = 4294967295; S = 6;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
#5 I0 = 4294967288; I1 = 4294967289; I2 = 4294967290; I3 = 4294967291; I4 = 4294967292; I5 = 4294967293; I6 = 4294967294; I7 = 4294967295; S = 7;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, S, Y);
end

endmodule