`timescale 1ns/1ps

module MUX32_32x1_TB;
wire [31:0] Y;
reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7;
reg [31:0] I8, I9, I10, I11, I12, I13, I14, I15;
reg [31:0] I16, I17, I18, I19, I20, I21, I22, I23;
reg [31:0] I24, I25, I26, I27, I28, I29, I30, I31;
reg [4:0] S;

MUX32_32x1 mux32_32x1_inst(.Y(Y), .I0(I0), .I1(I1), .I2(I2), .I3(I3),
                           .I4(I4), .I5(I5), .I6(I6), .I7(I7),
                           .I8(I8), .I9(I9), .I10(I10), .I11(I11),
                           .I12(I12), .I13(I13), .I14(I14), .I15(I15),
                           .I16(I16), .I17(I17), .I18(I18), .I19(I19),
                           .I20(I20), .I21(I21), .I22(I22), .I23(I23),
                           .I24(I24), .I25(I25), .I26(I26), .I27(I27),
                           .I28(I28), .I29(I29), .I30(I30), .I31(I31), .S(S));

initial
begin
I0 = 0; I1 = 0; I2 = 0; I3 = 0; I4 = 0; I5 = 0; I6 = 0; I7 = 0; I8 = 0; I9 = 0; I10 = 0; I11 = 0; I12 = 0; I13 = 0; I14 = 0; I15 = 0; I16 = 0; I17 = 0; I18 = 0; I19 = 0; I20 = 0; I21 = 0; I22 = 0; I23 = 0; I24 = 0; I25 = 0; I26 = 0; I27 = 0; I28 = 0; I29 = 0; I30 = 0; I31 = 0; S = 0;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 0;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 1;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 2;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 3;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 4;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 5;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 6;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 7;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 8;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 9;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 10;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 11;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 12;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 13;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 14;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 15;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 16;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 17;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 18;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 19;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 20;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 21;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 22;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 23;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 24;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 25;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 26;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 27;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 28;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 29;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 30;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
#5 I0 = 4294967264; I1 = 4294967265; I2 = 4294967266; I3 = 4294967267; I4 = 4294967268; I5 = 4294967269; I6 = 4294967270; I7 = 4294967271; I8 = 4294967272; I9 = 4294967273; I10 = 4294967274; I11 = 4294967275; I12 = 4294967276; I13 = 4294967277; I14 = 4294967278; I15 = 4294967279; I16 = 4294967280; I17 = 4294967281; I18 = 4294967282; I19 = 4294967283; I20 = 4294967284; I21 = 4294967285; I22 = 4294967286; I23 = 4294967287; I24 = 4294967288; I25 = 4294967289; I26 = 4294967290; I27 = 4294967291; I28 = 4294967292; I29 = 4294967293; I30 = 4294967294; I31 = 4294967295; S = 31;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d I16:%d I17:%d I18:%d I19:%d I20:%d I21:%d I22:%d I23:%d I24:%d I25:%d I26:%d I27:%d I28:%d I29:%d I30:%d I31:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
end

endmodule