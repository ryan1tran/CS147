`timescale 1ns/1ps

module MUX32_16x1_TB;
wire [31:0] Y;
reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7;
reg [31:0] I8, I9, I10, I11, I12, I13, I14, I15;
reg [3:0] S;

MUX32_16x1 mux32_16x1_inst(.Y(Y), .I0(I0), .I1(I1), .I2(I2), .I3(I3),
                           .I4(I4), .I5(I5), .I6(I6), .I7(I7),
                           .I8(I8), .I9(I9), .I10(I10), .I11(I11),
                           .I12(I12), .I13(I13), .I14(I14), .I15(I15), .S(S));

initial
begin
I0 = 0; I1 = 0; I2 = 0; I3 = 0; I4 = 0; I5 = 0; I6 = 0; I7 = 0; I8 = 0; I9 = 0; I10 = 0; I11 = 0; I12 = 0; I13 = 0; I14 = 0; I15 = 0; S = 0;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 0;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 1;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 2;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 3;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 4;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 5;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 6;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 7;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 8;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 9;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 10;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 11;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 12;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 13;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 14;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
#5 I0 = 4294967280; I1 = 4294967281; I2 = 4294967282; I3 = 4294967283; I4 = 4294967284; I5 = 4294967285; I6 = 4294967286; I7 = 4294967287; I8 = 4294967288; I9 = 4294967289; I10 = 4294967290; I11 = 4294967291; I12 = 4294967292; I13 = 4294967293; I14 = 4294967294; I15 = 4294967295; S = 15;
#5 $write("I0:%d I1:%d I2:%d I3:%d I4:%d I5:%d I6:%d I7:%d I8:%d I9:%d I10:%d I11:%d I12:%d I13:%d I14:%d I15:%d S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
end

endmodule