`timescale 1ns/1ps
// Name: mux32_16x1_tb.v
// Module: MUX32_16x1_TB
// Input: 
// Output: 
//
// Notes: Common definitions
// 
//
// Revision History:
//
// Version	Date		Who		email			note
//------------------------------------------------------------------------------------------
//  1.0     Apr 18, 2020	Ryan Tran	tranryanp@gmail.com	Initial creation
//------------------------------------------------------------------------------------------

module MUX32_16x1_TB;
reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15;
reg [3:0] S;
wire [31:0] Y;

MUX32_16x1 mux32_8x1_inst1(.Y(Y), .I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .I6(I6), .I7(I7), .I8(I8),
			   .I9(I9), .I10(I10), .I11(I11), .I12(I12), .I13(I13), .I14(I14), .I15(I15), .S(S));

initial
begin
I0 = 0; I1 = 0; I2 = 0; I3 = 0; I4 = 0; I5 = 0; I6 = 0; I7 = 0; I8 = 0; I9 = 0; I10 = 0; I11 = 0; I12 = 0; I13 = 0; I14 = 0; I15 = 0; S = 0;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 0;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 1;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 2;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 3;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 4;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 5;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 6;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 7;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 8;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 9;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 10;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 11;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 12;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 13;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 14;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; S = 15;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, S, Y);
end

endmodule
