`timescale 1ns/1ps
// Name: mux32_32x1_tb.v
// Module: MUX32_32x1_TB
// Input: 
// Output: 
//
// Notes: Common definitions
// 
//
// Revision History:
//
// Version	Date		Who		email			note
//------------------------------------------------------------------------------------------
//  1.0     Apr 18, 2020	Ryan Tran	tranryanp@gmail.com	Initial creation
//------------------------------------------------------------------------------------------

module MUX32_32x1_TB;
reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31;
reg [4:0] S;
wire [31:0] Y;

MUX32_32x1 mux32_32x1_inst1(.Y(Y), .I0(I0), .I1(I1), .I2(I2), .I3(I3),
                           .I4(I4), .I5(I5), .I6(I6), .I7(I7), .I8(I8),
			   .I9(I9), .I10(I10), .I11(I11), .I12(I12),
			   .I13(I13), .I14(I14), .I15(I15), .I16(I16),
			   .I17(I17), .I18(I18), .I19(I19), .I20(I20),
			   .I21(I21), .I22(I22), .I23(I23), .I24(I24),
			   .I25(I25), .I26(I26), .I27(I27), .I28(I28),
			   .I29(I29), .I30(I30), .I31(I31), .S(S));

initial
begin
I0 = 0; I1 = 0; I2 = 0; I3 = 0; I4 = 0; I5 = 0; I6 = 0; I7 = 0; I8 = 0; I9 = 0; I10 = 0; I11 = 0; I12 = 0; I13 = 0; I14 = 0; I15 = 0; I16 = 0; I17 = 0; I18 = 0; I19 = 0; I20 = 0; I21 = 0; I22 = 0; I23 = 0; I24 = 0; I25 = 0; I26 = 0; I27 = 0; I28 = 0; I29 = 0; I30 = 0; I31 = 0; S = 0;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 0;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 1;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 2;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 3;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 4;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 5;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 6;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 7;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 8;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 9;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 10;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 11;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 12;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 13;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 14;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 15;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 16;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 17;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 18;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 19;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 20;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 21;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 22;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 23;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 24;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 25;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 26;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 27;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 28;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 29;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 30;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
I0 = 1431655700; I1 = 1431655701; I2 = 1431655702; I3 = 1431655703; I4 = 1431655704; I5 = 1431655705; I6 = 1431655706; I7 = 1431655707; I8 = 1431655708; I9 = 1431655709; I10 = 1431655710; I11 = 1431655711; I12 = 1431655712; I13 = 1431655713; I14 = 1431655714; I15 = 1431655715; I16 = 1431655716; I17 = 1431655717; I18 = 1431655718; I19 = 1431655719; I20 = 1431655720; I21 = 1431655721; I22 = 1431655722; I23 = 1431655723; I24 = 1431655724; I25 = 1431655725; I26 = 1431655726; I27 = 1431655727; I28 = 1431655728; I29 = 1431655729; I30 = 1431655730; I31 = 1431655731; S = 31;
#5 $write("I0:%d, I1:%d, I2:%d, I3:%d, I4:%d, I5:%d, I6:%d, I7:%d, I8:%d, I9:%d, I10:%d, I11:%d, I12:%d, I13:%d, I14:%d, I15:%d, I16:%d, I17:%d, I17:%d, I18:%d, I20:%d, I21:%d, I22:%d, I23:%d, I24:%d, I25:%d, I26:%d, I27:%d, I28:%d, I29:%d, I30:%d, I31:%d, S:%d Y:%d\n", I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, S, Y);
end

endmodule
